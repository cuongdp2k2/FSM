module top (
    // input
    input logic clk_i ,
    input logic w_i   ,
    input logic res_ni ,

    // output
    output reg         z_o ,
    output reg [8:0] Stage_o 
);
	ex1 dut(
		.*
	);
	 
endmodule : top
