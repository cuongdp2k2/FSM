module top (
    // input
    input logic clk_i ,
    input logic w   ,
    input logic res_ni ,

    // output
    output reg         z_o ,
    output reg [3:0] State_o 
);
	ex2 dut(
		.*
	);
	 
endmodule : top
